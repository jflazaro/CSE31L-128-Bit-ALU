`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/29/2016 03:05:47 PM
// Design Name: 
// Module Name: FlagGen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FlagGen(
    input logic [2:0] opsel,
    input logic mode,
    input logic cin,
    output logic c_flag,
    output logic z_flag,
    output logic s_flag,
    output logic o_flag
    );
    
    
    
endmodule
